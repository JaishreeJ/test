module and_data(input a,input b,output c);
assign c = a & b;
endmodule
