module buffer_assign(input d,input enable,output y);
assign y=d;
endmodule
