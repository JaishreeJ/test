module andg_3(input a,input b,output c);
and x(c,a,b);
endmodule
