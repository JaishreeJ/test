module buffer1(input d,input enable,output y);
buf b1(y,enable,d);
endmodule
